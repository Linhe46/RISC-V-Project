/home/syetos/RISCV-Project/RTL/Common/mem.sv