/home/syetos/RISCV-Project/RTL/Common/registers.sv