/home/syetos/RISCV-Project/RTL/Common/wb.sv