/home/syetos/RISCV-Project/RTL/Common/id.sv