/home/syetos/RISCV-Project/RTL/Unique/RISCV-Trace/myCPU.sv