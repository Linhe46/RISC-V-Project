/home/syetos/RISCV-Project/RTL/Unique/RISCV-Trace/miniRV_SoC.sv