/home/syetos/RISCV-Project/RTL/Common/ex.sv