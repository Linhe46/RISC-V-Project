/home/syetos/RISCV-Project/RTL/Common/stall_unit.sv