/home/syetos/RISCV-Project/RTL/Unique/RISCV-Trace/mem_wb_reg.sv