/home/syetos/RISCV-Project/RTL/Unique/RISCV-Trace/ex_mem_reg.sv