/home/syetos/RISCV-Project/RTL/Common/forward_unit.sv