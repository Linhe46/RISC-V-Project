/home/syetos/RISCV-Project/RTL/Unique/RISCV-Trace/if_id_reg.sv