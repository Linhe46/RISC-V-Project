/home/syetos/RISCV-Project/RTL/Common/pc.sv