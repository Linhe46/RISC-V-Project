/home/syetos/RISCV-Project/RTL/Unique/RISCV-Trace/id_ex_reg.sv