/home/syetos/RISCV-Project/RTL/Common/bpd.sv